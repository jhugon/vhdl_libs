library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library neorv32;
use neorv32.neorv32_package.all;

entity neorv32_test_setup_bootloader is
  generic (
    -- adapt these for your setup --
    CLOCK_FREQUENCY   : natural := 100000000; -- clock frequency of clk_i in Hz
    MEM_INT_IMEM_SIZE : natural := 16*1024;   -- size of processor-internal instruction memory in bytes
    MEM_INT_DMEM_SIZE : natural := 8*1024     -- size of processor-internal data memory in bytes
  );
  port (
    -- Global control --
    clk       : in  std_ulogic; -- global clock, rising edge
    rstn_i      : in  std_ulogic; -- global reset, low-active, async
    sw : in std_ulogic_vector(15 downto 1); -- notice 0 is missing (it's rstn_i)
    -- GPIO --
    led      : out std_ulogic_vector(15 downto 0); -- parallel output
    -- UART0 --
    RsTx : out std_ulogic; -- UART0 send data
    RsRx : in  std_ulogic; -- UART0 receive data
    -- UART1 --
    UART1_tx : out std_ulogic;
    UART1_rx : in  std_ulogic
  );
end entity;

architecture neorv32_test_setup_bootloader_rtl of neorv32_test_setup_bootloader is

  signal con_gpio_i : std_ulogic_vector(63 downto 0);
  signal con_gpio_o : std_ulogic_vector(63 downto 0);

begin

  neorv32_top_inst: neorv32_top
  generic map (
    -- General --
    CLOCK_FREQUENCY              => CLOCK_FREQUENCY,   -- clock frequency of clk_i in Hz
    INT_BOOTLOADER_EN            => true,              -- boot configuration: true = boot explicit bootloader; false = boot from int/ext (I)MEM
    -- RISC-V CPU Extensions --
    CPU_EXTENSION_RISCV_C        => true,              -- implement compressed extension?
    CPU_EXTENSION_RISCV_M        => true,              -- implement mul/div extension?
    CPU_EXTENSION_RISCV_Zicsr    => true,              -- implement CSR system?
    CPU_EXTENSION_RISCV_Zicntr   => true,              -- implement base counters?
    -- Internal Instruction memory --
    MEM_INT_IMEM_EN              => true,              -- implement processor-internal instruction memory
    MEM_INT_IMEM_SIZE            => MEM_INT_IMEM_SIZE, -- size of processor-internal instruction memory in bytes
    -- Internal Data memory --
    MEM_INT_DMEM_EN              => true,              -- implement processor-internal data memory
    MEM_INT_DMEM_SIZE            => MEM_INT_DMEM_SIZE, -- size of processor-internal data memory in bytes
    -- Processor peripherals --
    IO_GPIO_EN                   => true,              -- implement general purpose input/output port unit (GPIO)?
    IO_MTIME_EN                  => true,              -- implement machine system timer (MTIME)?
    IO_UART0_EN                  => true,              -- implement primary universal asynchronous receiver/transmitter (UART0)?
    IO_UART1_EN                  => true,              -- implement primary universal asynchronous receiver/transmitter (UART1)?
    IO_UART1_RX_FIFO             => 8,                 -- add some extra to the fifo so that we don't need interrupts
    IO_UART1_TX_FIFO             => 8                  -- add some extra to the fifo so that we don't need interrupts
  )
  port map (
    -- Global control --
    clk_i       => clk,       -- global clock, rising edge
    rstn_i      => rstn_i,      -- global reset, low-active, async
    -- GPIO (available if IO_GPIO_EN = true) --
    gpio_i      => con_gpio_i,  -- parallel input
    gpio_o      => con_gpio_o,  -- parallel output
    -- primary UART0 (available if IO_UART0_EN = true) --
    uart0_txd_o => RsTx, -- UART0 send data
    uart0_rxd_i => RsRx, -- UART0 receive data
    uart1_txd_o => UART1_tx, -- UART1 send data
    uart1_rxd_i => UART1_rx  -- UART1 receive data
  );

  -- GPIO output --
  led <= con_gpio_o(15 downto 0);
  con_gpio_i <= "0000000000000000" & sw & '0' & con_gpio_o(31 downto 0);

end architecture;
